/home/ecegrid/a/mg106/ece337/Lab2/source/adder_nbit.sv